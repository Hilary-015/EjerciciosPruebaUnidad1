----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:48:41 05/23/2022 
-- Design Name: 
-- Module Name:    entidadPromedio2 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity entidadPromedio2 is
    Port ( A : in  STD_LOGIC_VECTOR (0 to 3);
           B : in  STD_LOGIC_VECTOR (0 to 3);
           C : out  STD_LOGIC_VECTOR (0 to 3));
end entidadPromedio2;

architecture Behavioral of entidadPromedio2 is

begin


end Behavioral;

