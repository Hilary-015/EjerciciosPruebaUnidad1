----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:46:14 05/23/2022 
-- Design Name: 
-- Module Name:    entidadProyecto - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity entidadProyecto is
    Port ( P0 : in  STD_LOGIC;
           P1 : in  STD_LOGIC;
           P2 : in  STD_LOGIC;
           A0 : out  STD_LOGIC;
           A1 : out  STD_LOGIC;
           X : inout  STD_LOGIC);
end entidadProyecto;

architecture Behavioral of entidadProyecto is

begin


end Behavioral;

